library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


entity corrector_1 is    
 port(    x : in std_logic_vector(0 to 15);
          c : in std_logic_vector(0 to 6);
          s : inout std_logic_vector(0 to 6);
          y : out std_logic_vector(0 to 15)    
     );      
end corrector_1;

architecture beh of corrector_1 is
    
    constant i0:std_logic_vector(0 to 6):="1000000";
    constant i1:std_logic_vector(0 to 6):="0100000";
    constant i2:std_logic_vector(0 to 6):="0010000";
    constant i3:std_logic_vector(0 to 6):="0001000";
    constant i4:std_logic_vector(0 to 6):="0000100";
    constant i5:std_logic_vector(0 to 6):="0000010";
    constant i6:std_logic_vector(0 to 6):="0000001";
   

  type par_chk_mat is array  (0 to 6) of std_logic_vector(0 to 22);
  signal h : par_chk_mat:=("10000001000100110011100",
                           "01000000101010101110010",
                           "00100001010001101001011",
                           "00010000100100011001000",
                           "00001001001100100001101",
                           "00000100110010001101010",
                           "00000010011001010110101");
  
  
  
    
 type look_up_table is array  (0 to 127) of std_logic_vector(0 to 15);
 signal l : look_up_table:=("0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
                            "0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000001100","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
                            "0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
                            "0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0011000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
                            "0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
                            "0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000",
                            "0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000001100000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000110000000000","0000000000000000",
                            "0000000000000000","0000000000000000","0000000000000000","0000000011000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","0000000000000000","1100000000000000","0000000000000000");
                            
   signal e : std_logic_vector(0 to 15);
 
      
begin

process(x,c,s,e)   
begin
 
  s(0)<=(((((((x(0) xor x(4)) xor x(7)) xor x(8)) xor x(11)) xor x(12)) xor x(13)) xor c(0));
  s(1)<=((((((((x(1) xor x(3)) xor x(5)) xor x(7)) xor x(9)) xor x(10)) xor x(11)) xor x(14)) xor c(1));
  s(2)<=((((((((x(0) xor x(2)) xor x(6)) xor x(7)) xor x(9)) xor x(12)) xor x(14)) xor x(15)) xor c(2));
  s(3)<=(((((x(1) xor x(4)) xor x(8)) xor x(9)) xor x(12)) xor c(3));
  s(4)<=(((((((x(0) xor x(3)) xor x(4)) xor x(7)) xor x(12)) xor x(13)) xor x(15)) xor c(4));
  s(5)<=(((((((x(1) xor x(2)) xor x(5)) xor x(9)) xor x(10)) xor x(12)) xor x(14)) xor c(5));
  s(6)<=((((((((x(2) xor x(3)) xor x(6)) xor x(8)) xor x(10)) xor x(11)) xor x(13)) xor x(15)) xor c(6));
  
  
  
  e<=l(conv_integer(s));
  
  y<=x  xor e;
   
      
end process;
  
end beh;
  

             
